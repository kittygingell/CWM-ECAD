//////////////////////////////////////////////////////////////////////////////////
// Exercise #2 - Doorbell Chime
// Student Name:
// Date: 
//
//  Description: In this exercise, you need to design a multiplexer that chooses between two sounds, where the  
//  output is delayed by 5 ticks (not clocks!) and acts according to the following truth table:
//
//  sel | out
// -----------------
//   0  | a
//   1  | b
//
//  inputs:
//           a, b, sel
//
//  outputs:
//           out
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

//Defining the module

module doorbell(
	input a,
	input b,
	input sel,
	output out);
 
//Registers and wires
  
	reg r;
	wire out;
	
//Logic
			always @(sel or a or b);
			begin
				if (sel == 1)
					r <= b;
				else
					r <= a;
			end

		assign #5 out=r;    
      
endmodule
